--Generic Register with synchronous reset

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity DATA_REGISTER is
	generic (data_width:integer);
	port(
			clk:	in std_logic;
			reset: 	in std_logic;
			enable: in std_logic;			
			Din: 	in std_logic_vector(data_width-1 downto 0);
			
	      	Dout: 	out std_logic_vector(data_width-1 downto 0)
	      	
	     );
end entity;


architecture Behave of DATA_REGISTER is
begin
	
	process(clk)
    begin
       if(clk'event and (clk  = '1')) then
       	   if(reset = '0') then
       	   		Dout <= std_logic_vector(to_unsigned(0,data_width));
       	   		
           elsif(enable = '1') then           
           		Dout <= Din;           		           
           end if;                      
       end if;          
    end process;
end Behave;

